    Mac OS X            	   2   �      �                                      ATTR D�5   �   �   -                  �   -  com.apple.quarantine q/0000;4be3e883;Safari.app;|com.apple.Safari 