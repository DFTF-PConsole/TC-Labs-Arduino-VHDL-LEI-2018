    Mac OS X            	   2   �      �                                      ATTR e,�   �   �   I                  �   I  com.apple.quarantine q/0000;506beff3;Mail;7D2E3DC3-0B34-4801-8F55-153E898F40AB|com.apple.mail 